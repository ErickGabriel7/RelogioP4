--Autor: Erick Gabriel
-- teste de leds
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY relogiop4 IS
PORT( CLOCK_50 : IN STD_LOGIC;
      KEY      : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      LEDR     : OUT STD_LOGIC_VECTOR(8 DOWNTO 0));

END relogiop4;

ARCHITECTURE imp OF relogiop4 IS
COMPONENT pll1m is
	port (
		refclk   : in  std_logic := '0'; --  refclk.clk
		rst      : in  std_logic := '0'; --   reset.reset
		outclk_0 : out std_logic;        -- outclk0.clk
		locked   : out std_logic         --  locked.export
	);
END COMPONENT;

COMPONENT div5b IS
PORT( rst,clk : IN  STD_LOGIC;
      q       : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
END COMPONENT;

SIGNAL RST50, RST : STD_LOGIC;
SIGNAL q1, q2, q3, q4  :  STD_LOGIC_VECTOR(4 DOWNTO 0);
SIGNAL contador        :  STD_LOGIC_VECTOR(19 DOWNTO 0);
SIGNAL clk             :  STD_LOGIC;
BEGIN
PROCESS(Clock_50)
   BEGIN
	  IF CLOCK_50'EVENT AND CLOCK_50 = '1' THEN
	    RST50 <= NOT KEY(0);
	  END IF;
	END PROCESS;
	
	PLL0 : pll1m PORT MAP (
	   refclk   => CLOCK_50,
		rst      => rst50,
		outclk_0 => clk,
		locked   => rst);
		
	 u0: div5b PORT MAP(rst => rst, clk => clk  , q => q1);
    u1: div5b PORT MAP(rst => rst, clk => q1(4), q => q2);
    u2: div5b PORT MAP(rst => rst, clk => q2(4), q => q3);
    u3: div5b PORT MAP(rst => rst, clk => q3(4), q => q4);
    contador <= q4 & q3 & q2 & q1;
	 LEDR <= contador(19 DOWNTO 11);
END imp;

